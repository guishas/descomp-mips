library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM IS
   generic (
          dataWidth: natural := 32;
          addrWidth: natural := 32;
			 memoryAddrWidth:  natural := 6 -- 64 posicoes de 32 bits cada 
	);   
   port (
          Endereco : in  std_logic_vector (addrWidth-1 downto 0);
          Dado     : out std_logic_vector (dataWidth-1 downto 0) 		 
	);
end entity;

architecture assincrona OF ROM IS
	type blocoMemoria IS ARRAY(0 TO 2**memoryAddrWidth - 1) OF std_logic_vector(dataWidth-1 downto 0);

	function initMemory
		return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
	begin

		tmp(0)  := "000000" & "00000" & "00000" & "00000" & "00000" & "000000"; -- NOP
		tmp(1)  := "000000" & "01011" & "01010" & "01001" & "00000" & "100000"; -- SOMA
		tmp(2)  := "000000" & "01011" & "01010" & "01001" & "00000" & "100010"; -- SUB
		tmp(3)  := "000000" & "00000" & "00000" & "00000" & "00000" & "000000"; -- NOP
		tmp(4)  := "000000" & "01011" & "01010" & "0000000001000000"; -- SW
		tmp(5)  := "000000" & "00000" & "00000" & "0000000000000000"; -- NOP
		tmp(6)  := "000000" & "01011" & "01010" & "0000000001000000"; -- LW
		tmp(7)  := "000000" & "01010" & "01010" & "0000000000000010"; -- BEQ
		tmp(10) := "000000" & "00000" & "00000" & "0000000000000000"; -- NOP
		tmp(11) := "000000" & "00000000000000000000000000"; -- J

		return tmp;
   end initMemory;


   signal memROM : blocoMemoria := initMemory;   
	signal EnderecoLocal : std_logic_vector(memoryAddrWidth-1 downto 0);

begin

  EnderecoLocal <= Endereco(memoryAddrWidth+1 downto 2);
  Dado <= memROM (to_integer(unsigned(EnderecoLocal)));
  
end architecture;
